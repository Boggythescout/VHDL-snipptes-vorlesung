architecture medwedew of puls is

begin
