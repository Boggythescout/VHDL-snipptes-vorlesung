entity puls is 
	port(
		clk, x, res_n: in std_logic;
		y: out std_logic
		);
end entity puls;

architecture medwedew of puls is
begin
	
