entity mux is 
	port(
		s, e0, e1, e2: in std_logic;
		a: out std_logic
		);
end entity mux;